library IEEE;
-- Please add necessary libraries:


entity controller is
    port (
        clk         : in    std_logic;
        reset       : in    std_logic;

        sensor_l    : in    std_logic;
        sensor_m    : in    std_logic;
        sensor_r    : in    std_logic;

        count_in    : in    std_logic_vector (?? downto 0);  -- Please enter upper bound
        count_reset : out   std_logic;

        motor_l_reset       : out   std_logic;
        motor_l_direction   : out   std_logic;

        motor_r_reset       : out   std_logic;
        motor_r_direction   : out   std_logic
    );
end entity controller;
